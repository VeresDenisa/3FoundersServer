package base_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "base_agent_config.svh"

  `include "base_driver.svh"
  `include "base_monitor.svh"
  
  `include "base_agent.svh"
endpackage : base_pack;