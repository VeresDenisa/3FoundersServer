package port_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "port_driver.svh"
  `include "port_monitor.svh"
  `include "port_sequencer.svh"

  `include "port_agent.svh"
endpackage : port_agent_pack;