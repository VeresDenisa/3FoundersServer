package item_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "src/test/item/data_packet.svh"
  `include "src/test/item/control_item.svh"
  `include "src/test/item/memory_item.svh"
  `include "src/test/item/reset_item.svh"
  `include "src/test/item/port_item.svh"
endpackage : item_pack;