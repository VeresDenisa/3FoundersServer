package memory_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "memory_driver.svh"
  `include "memory_monitor.svh"

  `include "memory_agent.svh"
endpackage : memory_agent_pack;