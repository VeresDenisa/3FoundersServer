package reset_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "reset_driver.svh"
  `include "reset_monitor.svh"

  `include "reset_agent.svh"
endpackage : reset_agent_pack;