package env_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import seq_pack::*;
  import base_pack::*;
  import config_pack::*;

  import reset_agent_pack::*;
  import control_agent_pack::*;
  import memory_agent_pack::*;
  import port_agent_pack::*;

  `include "virtual_sequencer.svh"
  `include "virtual_sequence.svh"

  `include "scoreboard.svh"

  `include "port_covergroup.sv"
  `include "control_covergroup.sv"
  `include "memory_covergroup.sv"
  `include "data_covergroup.sv"
  `include "event_covergroup.sv" 

  `include "port_coverage.svh"
  `include "coverage.svh"

  `include "environment.svh"
endpackage : env_pack;