package control_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "control_driver.svh"
  `include "control_monitor.svh"

  `include "control_agent.svh"
endpackage : control_agent_pack;