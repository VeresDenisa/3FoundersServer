package memory_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "src/test/environment/agent_memory/memory_driver.svh"
  `include "src/test/environment/agent_memory/memory_monitor.svh"

  `include "src/test/environment/agent_memory/memory_agent.svh"
endpackage : memory_agent_pack;