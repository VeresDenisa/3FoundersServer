package item_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "data_packet.svh"
  `include "control_item.svh"
  `include "memory_item.svh"
  `include "reset_item.svh"
  `include "port_item.svh"
endpackage : item_pack;